module config_reg(
    input  Logic clk,
    input  Logic reset,
    input  Logic write,
    input  Logic [15:0] data_in,
    input  Logic [2:0] address,
    output Logic [15:0] data_out
);

protected

MTTI;HDU;Wt?N\Ev)p$.,h.Rg#"cok2*.fUl '?K9?"kDn2YBkJWI,k7+DJ.[a92?\Tko^#4"m1t^VEU
Y-,Jeo-mnc;onWIzUp!k$>TBlVIA6ba9Ia??],5XuOkyL77P?1aeksKoz[,vCYV5WCABAKE=5QA@
!dsa]#l+1r+pvrAZeEgwAqLD\EXU7fV5+I4t+B-kkX-+KXvWov)[0d]JuJv2c96,I(1J,DZ$74,o
C!q?[_Xpe_KwGpw4EaAlRT3S3sti_Si.rv17*RY8kXeV0W2xm]!adglo2L!J2"d~]Vy;%&*Y
?+nA?Iell1ZP1"+rrT=1ekstP+O;JpaM,.sz,V02!_l3eby$jrsih~%QTp-lle^X$"2}EVT!
??_ab.a1'^z7AKR2nb;.Voo^P+vz2MDU;SrIanI mI"J0~ hslo"ei;v07WL9CwGnf;L"!ka#\
E2HI;yU2x5HaliVGj}{KE2wvJUzTHk3e62s0Jc5Q[BAuWlo?eeU3D2LtP(5NcEkNejt4??7
Z>2ZKp_"xK.Ki2Z2^2vv)5W#[;fwq2sA{twO FLX^WE3,>oo"JKVvW+.)9E~C2P!p)??0,
+b*#W+QASi ~8O%Rw9j,=]5?BRt4,wUhAW^x9xO5qZJXQ[0sbXBdw!P0w(,FgZXm(Az'\n~
r98jh2Hxo~.T$0hWnI{ny>M\Mf-=b!{}L??g2Uf1^J$l) y}{gJ5H)Zlpl0jX<]{6)+:
qk>M"I)9OXealLS8O>2YJ1Ti~U*99!ec4*(]/(l$ZN@?KPxPVrTHT_d!rsCJeX#Vl+C7(;
W??Y/!^rDs_n^urN@&Jc_1^mbU"UDt(=2^x?duE5z9+01DE3IP[+}7|p+TtO7)?2"7Wdbu.
zi3"^t5skv1NLteWSX <dZkeepY"[OwRVpkl*0qyF]!OjO0FsrOPJpC,mlrp*"4mpEt'4
1]@*L>!5K?;igVsu!n08y;TTW1c#9oAO2EZs;Wz0aQ*U0L?=DP5$H2~KQ?;,;t+]BA)*
<Epq:(!OH0pJpr"_=}pmSxZBHK",rCikEY)_lrF,}wrPCkQU)9~sB".g.2pa-DlI.Vu?0
nA:jzMwH}1yIcsaN!5r+21zPmT.bB1xYnoGVq,qAO2]E;[r.~D~5YAjsVJrssI?L\_M/H
3w0)K]Gs,Yo!+RE77XKG+"A5i7;KBo@q=i

endprotected

endmodule // test