///////////////////////////////////////////////////////////////////////////////
// Author: Kareem Waseem
// Course: Digital Verification using SV & UVM
//
// Description: Counter Design
///////////////////////////////////////////////////////////////////////////////

module counter (clk, rst_n, load_n, up_down, ce, data_load, count_out, max_count, zero);
parameter WIDTH = 4;

input clk;
input rst_n;
input load_n;
input up_down;
input ce;
input [WIDTH-1:0] data_load;
output reg [WIDTH-1:0] count_out;
output max_count;
output zero;

always @(posedge clk) begin
    if (!rst_n)
        count_out <= 0;
    else if (!load_n)
        count_out <= data_load;
    else if (ce) begin
        if (up_down)
            count_out <= count_out + 1;
        else
            count_out <= count_out - 1;
    end
end

assign max_count = (count_out == {WIDTH{1'b1}}) ? 1 : 0;
assign zero      = (count_out == 0) ? 1 : 0;

endmodule