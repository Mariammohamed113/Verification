package constant_enums;

typedef enum { OR, XOR, ADD, MULT, SHIFT, ROTATE, INVALID6, INVALID7 } Opcode_e;

typedef enum {MAXPOS=3, MAXNEG=-4, ZERO=0} corner_state_e;

endpackage